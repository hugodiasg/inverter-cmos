*INVERTER CMOS

.subckt inverter_post	IN	OUT	VCC	VGND	VSUBS

M1	OUT	IN	VCC	VCC	pshort_model	w=3u l=0.15u
M2	OUT	IN	VGND	VGND	nshort_model	w=1u l=0.15u

C0 IN VDD 0.03fF
C1 IN GND 0.02fF
C2 VDD OUT 0.29fF
C3 GND OUT 0.11fF
C4 IN OUT 0.05fF
C5 GND VSUBS 0.29fF
C6 OUT VSUBS 0.13fF
C7 VDD VSUBS 0.39fF
C8 IN VSUBS 0.30fF
*C9 w_n36_344# VSUBS 0.52fF
.ends
